`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/09/2023 10:28:02 AM
// Design Name: 
// Module Name: TopLevel_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module TopLevel_tb(
    );
    
    parameter n = 32;
    reg clk;
    reg [2:0] op;
    reg [n - 1 : 0] R2;
    reg [n - 1 : 0] R3;
    wire [n - 1 : 0] R0;
    
    wire [n - 1 : 0] ResultVerify;
    wire ErrorFlag;
    
    TopLevel top(.R0(R0), .R2(R2), .R3(R3), .op(op), .clk(clk));
    
    // Verification 
    Verification verify (.Result(ResultVerify), .clk(clk), .op(op), .R2(R2), .R3(R3));
    
    assign ErrorFlag = (R0 != ResultVerify);

    always @ (posedge clk) begin
        if (ErrorFlag)
            $display("Error occurs when op = %d, R2 = %d, R3 = %d", op, R2, R3);
        end
    
    initial begin
        /*
        R2 = 0; R3 = 0; clk = 0;
        op = 3'b010;
        #100 op = 3'b001;
        */
        R2 = 32'b0; R3 = 32'b0; op = 3'b000; clk = 1'b0;
        #25 R2 = 32'b11010000101000010000101011101010; 
        
        #25 op = 3'b001;
        R2 = 32'b11111111111111111111111111111111;

        #25 op = 3'b010;
        R2 = 32'b00111011100110101100101000000000; // 1,000,000,000
        R3 = 32'b00111011100110101100101000000000; // 1,000,000,000

        #25 R2 = 32'b01000000000000000000000000000000; //1,073,741,824
        R3 = 32'b01000000000000000000000000000000; //1,073,741,824

        #25 R2 = 32'b00000000000000000000000000001101; // 13
        R3 = 32'b00000000000000000000000000001111; // 15

        #25 R2 = 32'b11111111111111111111111110100000; //-96
        R3 = 32'b00000000000000000000000000011100; //28
        
        #25 op = 3'b011;
        R2 = 32'b01101010111101100000100101011111; //1,794,509,151
        R3 = 32'b01101010111101100000100101011111; //1,794,509,151

        #25 R2 = 32'b01101010111101100000100101011111; // 1,794,509,151
        R3 = 32'b01110001010010100110001010001100; // -1,900,700,300
    
        #25 R2 = 32'b01101010111101100000100101011111; //1,794,509,151
        R3 = 32'b01011111011010100001001001100000; //1,600,787,040

        #25 R2 = 32'b00000000000010101111011010101111;
        R3 = 32'b00000000000000000000000000000000;

        #25 op = 3'b100;
        R2 = 32'b01010000101011111000011010011100; // 1353680540
        R3 = 32'b00100001111110000000010101101001; // 569902441
     
        #25 op = 3'b101;
        R2 = 32'b01010010000011111001011010100101; 
        R3 = 32'b01010000101011111000011010011100;
  
    end
    
    always #3 clk = ~clk;
    
endmodule
